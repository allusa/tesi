//: version "1.8.7"

module disc4max(D1, consolida, D2, nouv, D3, valor, D0);
//: interface  /sz:(159, 169) /bd:[ Li0>consolida(144/169) Li1>nouv(66/169) Li2>valor[7:0](30/169) Ro0<D3[7:0](110/169) Ro1<D2[7:0](82/169) Ro2<D1[7:0](54/169) Ro3<D0[7:0](26/169) ]
input [7:0] valor;    //: /sn:0 {0}(-110,78)(-25,78){1}
//: {2}(-21,78)(30,78){3}
//: {4}(-23,76)(-23,26)(145,26)(145,32){5}
supply0 w15;    //: /sn:0 {0}(194,109)(209,109)(209,129){1}
output [7:0] D2;    //: /sn:0 /dp:1 {0}(385,275)(385,267){1}
//: {2}(387,265)(536,265)(536,266)(548,266){3}
//: {4}(385,263)(385,257){5}
output [7:0] D1;    //: /sn:0 /dp:1 {0}(385,236)(385,226){1}
//: {2}(387,224)(465,224)(465,222)(546,222){3}
//: {4}(385,222)(385,215){5}
supply0 w0;    //: /sn:0 {0}(440,314)(440,292){1}
//: {2}(440,288)(440,253){3}
//: {4}(440,249)(440,211){5}
//: {6}(440,207)(440,167)(424,167){7}
//: {8}(438,209)(424,209){9}
//: {10}(438,251)(424,251){11}
//: {12}(438,290)(424,290){13}
input nouv;    //: /sn:0 {0}(-111,104)(118,104){1}
output [7:0] D0;    //: /sn:0 /dp:1 {0}(385,194)(385,184){1}
//: {2}(387,182)(505,182)(505,181)(544,181){3}
//: {4}(385,180)(385,173){5}
input consolida;    //: /sn:0 {0}(-101,326)(281,326)(281,164){1}
//: {2}(283,162)(314,162)(314,162)(340,162){3}
//: {4}(344,162)(348,162){5}
//: {6}(342,164)(342,202){7}
//: {8}(344,204)(348,204){9}
//: {10}(342,206)(342,244){11}
//: {12}(344,246)(348,246){13}
//: {14}(342,248)(342,285)(348,285){15}
//: {16}(281,160)(281,99)(225,99){17}
output [7:0] D3;    //: /sn:0 /dp:1 {0}(548,315)(385,315)(385,296){1}
supply1 w2;    //: /sn:0 {0}(424,199)(450,199){1}
//: {2}(452,197)(452,159){3}
//: {4}(452,155)(452,137){5}
//: {6}(450,157)(424,157){7}
//: {8}(452,201)(452,239){9}
//: {10}(450,241)(424,241){11}
//: {12}(452,243)(452,280)(424,280){13}
wire [7:0] w14;    //: /sn:0 {0}(30,46)(14,46){1}
//: {2}(12,44)(12,5)(165,5)(165,32){3}
//: {4}(12,48)(12,145)(153,145){5}
//: {6}(157,145)(385,145)(385,152){7}
//: {8}(155,143)(155,115){9}
wire w23;    //: /sn:0 {0}(132,48)(86,48){1}
wire [7:0] w24;    //: /sn:0 {0}(155,61)(155,94){1}
wire w18;    //: /sn:0 {0}(96,77)(86,77){1}
wire w8;    //: /sn:0 {0}(209,99)(194,99){1}
//: enddecls

  //: supply1 g4 (w2) @(463,137) /sn:0 /w:[ 5 ]
  register g8 (.Q(D3), .D(D2), .EN(w0), .CLR(w2), .CK(consolida));   //: @(385,285) /sn:0 /w:[ 1 0 13 13 15 ]
  //: joint g13 (D1) @(385, 224) /w:[ 2 4 -1 1 ]
  //: joint g37 (w14) @(12, 46) /w:[ 1 2 -1 4 ]
  //: joint g34 (consolida) @(281, 162) /w:[ 2 16 -1 1 ]
  //: frame g2 @(-40,-32) /sn:0 /wi:279 /ht:227 /tx:""
  register g1 (.Q(D0), .D(w14), .EN(w0), .CLR(w2), .CK(consolida));   //: @(385,162) /sn:0 /w:[ 5 7 7 7 5 ]
  //: joint g16 (w2) @(452, 241) /w:[ -1 9 10 12 ]
  not g28 (.I(consolida), .Z(w8));   //: @(219,99) /sn:0 /R:2 /w:[ 17 0 ]
  register g32 (.Q(w14), .D(w24), .EN(w15), .CLR(w8), .CK(nouv));   //: @(155,104) /sn:0 /w:[ 9 1 0 1 1 ]
  //: comment g27 /dolink:0 /link:"" @(387,106) /sn:0
  //: /line:"Disc"
  //: /end
  //: joint g19 (w0) @(440, 251) /w:[ -1 4 10 3 ]
  //: output g38 (D1) @(543,222) /sn:0 /w:[ 3 ]
  register g6 (.Q(D1), .D(D0), .EN(w0), .CLR(w2), .CK(consolida));   //: @(385,204) /sn:0 /w:[ 5 0 9 0 9 ]
  //: joint g9 (D0) @(385, 182) /w:[ 2 4 -1 1 ]
  register g7 (.Q(D2), .D(D1), .EN(w0), .CLR(w2), .CK(consolida));   //: @(385,246) /sn:0 /w:[ 5 0 11 11 13 ]
  //: input g31 (consolida) @(-103,326) /sn:0 /w:[ 0 ]
  //: joint g20 (w0) @(440, 209) /w:[ -1 6 8 5 ]
  //: joint g15 (w2) @(452, 199) /w:[ -1 2 1 8 ]
  //: comment g39 /dolink:0 /link:"" @(194,-60) /sn:0
  //: /line:"Disc atribut"
  //: /end
  //: output g43 (D2) @(545,266) /sn:0 /w:[ 3 ]
  //: input g25 (nouv) @(-113,104) /sn:0 /w:[ 0 ]
  //: supply0 g17 (w0) @(440,320) /sn:0 /w:[ 0 ]
  //: comment g29 /dolink:0 /link:"" @(78,-27) /sn:0
  //: /line:"Buffer"
  //: /end
  //: joint g42 (valor) @(-23, 78) /w:[ 2 4 1 -1 ]
  //: joint g5 (w2) @(452, 157) /w:[ -1 4 6 3 ]
  //: joint g14 (D2) @(385, 265) /w:[ 2 4 -1 1 ]
  //: output g44 (D3) @(545,315) /sn:0 /w:[ 0 ]
  //: input g24 (valor) @(-112,78) /sn:0 /w:[ 0 ]
  //: frame g36 @(-73,-65) /sn:0 /wi:574 /ht:450 /tx:""
  //: joint g21 (consolida) @(342, 204) /w:[ 8 7 -1 10 ]
  //: supply0 g23 (w15) @(209,135) /sn:0 /w:[ 1 ]
  //: joint g41 (w14) @(155, 145) /w:[ 6 8 5 -1 ]
  //: comment g40 /dolink:0 /link:"" @(78,-14) /sn:0
  //: /line:"Màxim"
  //: /end
  //: output g0 (D0) @(541,181) /sn:0 /w:[ 3 ]
  //: frame g26 @(328,104) /sn:0 /wi:158 /ht:235 /tx:""
  //: joint g22 (consolida) @(342, 246) /w:[ 12 11 -1 14 ]
  mux g35 (.I0(valor), .I1(w14), .S(w23), .Z(w24));   //: @(155,48) /sn:0 /w:[ 5 3 0 0 ] /ss:0 /do:0
  //: joint g18 (w0) @(440, 290) /w:[ -1 2 12 1 ]
  //: joint g30 (consolida) @(342, 162) /w:[ 4 -1 3 6 ]
  CMP8 g33 (.A(w14), .B(valor), .AgB(w23), .AeqB(w18));   //: @(31, 34) /sz:(54, 60) /sn:0 /p:[ Li0>0 Li1>3 Ro0<1 Ro1<1 ]

endmodule

module CMP8(AeqB, AgB, B, A);
//: interface  /sz:(54, 60) /bd:[ Li0>A[7:0](12/60) Li1>B[7:0](44/60) Ro0<AgB(14/60) Ro1<AeqB(43/60) ]
input [7:0] B;    //: /sn:0 {0}(100,142)(146,142)(146,211){1}
//: {2}(146,212)(146,333){3}
//: {4}(146,334)(146,387){5}
input [7:0] A;    //: /sn:0 /dp:2 {0}(99,115)(119,115)(119,175){1}
//: {2}(119,176)(119,239)(118,239)(118,300){3}
//: {4}(118,301)(118,378){5}
output AeqB;    //: /sn:0 {0}(527,407)(432,407){1}
output AgB;    //: /sn:0 {0}(530,370)(418,370)(418,363){1}
wire w6;    //: /sn:0 /dp:1 {0}(411,409)(302,409)(302,326)(292,326){1}
wire [3:0] w4;    //: /sn:0 {0}(122,301)(130,301)(130,297)(220,297){1}
wire [3:0] w0;    //: /sn:0 {0}(123,176)(221,176){1}
wire [3:0] w1;    //: /sn:0 {0}(150,212)(221,212){1}
wire w8;    //: /sn:0 {0}(293,174)(408,174)(408,334){1}
wire w2;    //: /sn:0 {0}(428,334)(428,295)(292,295){1}
wire w13;    //: /sn:0 /dp:1 {0}(395,350)(342,350){1}
//: {2}(340,348)(340,205)(293,205){3}
//: {4}(340,352)(340,404)(411,404){5}
wire [3:0] w5;    //: /sn:0 {0}(150,334)(158,334)(158,333)(220,333){1}
//: enddecls

  A4CMPB4 g4 (.B(w1), .A(w0), .AeqB(w13), .AgB(w8));   //: @(222, 162) /sz:(70, 65) /sn:0 /p:[ Li0>1 Li1>1 Ro0<3 Ro1<0 ]
  tran g8(.Z(w4), .I(A[3:0]));   //: @(116,301) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: output g3 (AeqB) @(524,407) /sn:0 /w:[ 0 ]
  mux g13 (.I0(w8), .I1(w2), .S(w13), .Z(AgB));   //: @(418,350) /sn:0 /w:[ 1 0 0 1 ] /ss:0 /do:0
  //: output g2 (AgB) @(527,370) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(98,142) /sn:0 /w:[ 0 ]
  //: joint g11 (w13) @(340, 350) /w:[ 1 2 -1 4 ]
  and g10 (.I0(w13), .I1(w6), .Z(AeqB));   //: @(422,407) /sn:0 /w:[ 5 0 1 ]
  tran g6(.Z(w1), .I(B[7:4]));   //: @(144,212) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  A4CMPB4 g7 (.B(w5), .A(w4), .AeqB(w6), .AgB(w2));   //: @(221, 283) /sz:(70, 65) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<1 ]
  tran g9(.Z(w5), .I(B[3:0]));   //: @(144,334) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  tran g5(.Z(w0), .I(A[7:4]));   //: @(117,176) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: input g0 (A) @(97,115) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire [7:0] w6;    //: /sn:0 {0}(492,166)(492,178)(467,178)(467,136)(295,136){1}
wire w7;    //: /sn:0 {0}(131,415)(21,415){1}
wire [7:0] w16;    //: /sn:0 {0}(489,426)(489,435)(458,435)(458,382)(292,382){1}
wire [7:0] w15;    //: /sn:0 {0}(492,333)(492,343)(466,343)(466,325)(292,325){1}
wire [7:0] w4;    //: /sn:0 {0}(495,75)(495,80)(295,80){1}
wire [7:0] w3;    //: /sn:0 {0}(494,115)(494,129)(468,129)(468,108)(295,108){1}
wire w0;    //: /sn:0 {0}(42,120)(134,120){1}
wire [7:0] w1;    //: /sn:0 {0}(491,288)(491,297)(292,297){1}
wire [7:0] w8;    //: /sn:0 {0}(491,378)(491,388)(466,388)(466,353)(292,353){1}
wire w2;    //: /sn:0 {0}(39,198)(60,198){1}
//: {2}(64,198)(134,198){3}
//: {4}(62,200)(62,337)(131,337){5}
wire [7:0] w10;    //: /sn:0 {0}(20,74)(20,84)(134,84){1}
wire w5;    //: /sn:0 {0}(-120,-29)(-44,-29)(-44,-41){1}
wire [7:0] w9;    //: /sn:0 /dp:1 {0}(492,216)(492,228)(461,228)(461,164)(350,164){1}
//: {2}(346,164)(295,164){3}
//: {4}(348,166)(348,247)(92,247)(92,301)(131,301){5}
//: enddecls

  led g8 (.I(w15));   //: @(492,326) /sn:0 /w:[ 0 ] /type:2
  //: joint g4 (w2) @(62, 198) /w:[ 2 -1 1 4 ]
  led g3 (.I(w4));   //: @(495,68) /sn:0 /w:[ 0 ] /type:2
  //: joint g2 (w9) @(348, 164) /w:[ 1 -1 2 4 ]
  disc4max g1 (.valor(w9), .nouv(w2), .consolida(w7), .D0(w1), .D1(w15), .D2(w8), .D3(w16));   //: @(132, 271) /sz:(159, 169) /sn:0 /p:[ Li0>5 Li1>5 Li2>0 Ro0<1 Ro1<1 Ro2<1 Ro3<1 ]
  led g11 (.I(w6));   //: @(492,159) /sn:0 /w:[ 0 ] /type:2
  led g10 (.I(w3));   //: @(494,108) /sn:0 /w:[ 0 ] /type:2
  led g6 (.I(w1));   //: @(491,281) /sn:0 /w:[ 0 ] /type:2
  //: dip g38 (w10) @(20,64) /sn:0 /w:[ 0 ] /st:2
  led g9 (.I(w16));   //: @(489,419) /sn:0 /w:[ 0 ] /type:2
  led g7 (.I(w8));   //: @(491,371) /sn:0 /w:[ 0 ] /type:2
  //: switch g31 (w0) @(25,120) /sn:0 /w:[ 0 ] /st:0
  disc4max g43 (.valor(w10), .nouv(w0), .consolida(w2), .D0(w4), .D1(w3), .D2(w6), .D3(w9));   //: @(135, 54) /sz:(159, 169) /sn:0 /p:[ Li0>1 Li1>1 Li2>3 Ro0<1 Ro1<1 Ro2<1 Ro3<3 ]
  led g25 (.I(w5));   //: @(-44,-48) /sn:0 /w:[ 1 ] /type:0
  //: switch g5 (w7) @(4,415) /sn:0 /w:[ 1 ] /st:0
  clock g24 (.Z(w5));   //: @(-133,-29) /sn:0 /w:[ 0 ] /omega:1000 /phi:0 /duty:50
  //: switch g0 (w2) @(22,198) /sn:0 /w:[ 0 ] /st:0
  led g12 (.I(w9));   //: @(492,209) /sn:0 /w:[ 0 ] /type:2

endmodule

module A4CMPB4(AgB, B, AeqB, A);
//: interface  /sz:(70, 65) /bd:[ Li0>B[3:0](50/65) Li1>A[3:0](14/65) Ro0<AeqB(43/65) Ro1<AgB(12/65) ]
input [3:0] B;    //: /sn:0 {0}(88,76)(157,76)(157,100){1}
//: {2}(157,101)(157,125){3}
//: {4}(157,126)(157,151){5}
//: {6}(157,152)(157,178){7}
//: {8}(157,179)(157,229){9}
//: {10}(157,230)(157,253){11}
//: {12}(157,254)(157,277){13}
//: {14}(157,278)(157,299){15}
//: {16}(157,300)(157,318){17}
input [3:0] A;    //: /sn:0 {0}(88,46)(123,46)(123,95){1}
//: {2}(123,96)(123,120){3}
//: {4}(123,121)(123,146){5}
//: {6}(123,147)(123,173){7}
//: {8}(123,174)(123,223){9}
//: {10}(123,224)(123,245){11}
//: {12}(123,246)(123,271){13}
//: {14}(123,272)(123,295){15}
//: {16}(123,296)(123,313){17}
output AeqB;    //: /sn:0 {0}(614,275)(537,275){1}
output AgB;    //: /sn:0 /dp:1 {0}(481,107)(607,107){1}
wire w32;    //: /sn:0 {0}(367,156)(391,156)(391,106)(411,106){1}
wire w6;    //: /sn:0 {0}(161,126)(186,126){1}
wire w7;    //: /sn:0 {0}(127,147)(225,147){1}
wire w16;    //: /sn:0 {0}(246,276)(382,276){1}
//: {2}(386,276)(414,276){3}
//: {4}(384,274)(384,188)(396,188){5}
wire w14;    //: /sn:0 {0}(127,272)(171,272)(171,273)(225,273){1}
wire w4;    //: /sn:0 /dp:1 {0}(295,124)(246,124){1}
wire w15;    //: /sn:0 {0}(161,278)(225,278){1}
wire w38;    //: /sn:0 /dp:1 {0}(225,126)(202,126){1}
wire w3;    //: /sn:0 /dp:1 {0}(161,101)(187,101){1}
wire w37;    //: /sn:0 /dp:1 {0}(414,281)(311,281)(311,299)(245,299){1}
wire w34;    //: /sn:0 {0}(204,152)(225,152){1}
wire w21;    //: /sn:0 /dp:1 {0}(346,153)(316,153){1}
wire w31;    //: /sn:0 /dp:1 {0}(396,183)(368,183){1}
wire w28;    //: /sn:0 {0}(295,182)(275,182){1}
//: {2}(273,180)(273,157){3}
//: {4}(275,155)(295,155){5}
//: {6}(273,153)(273,129)(295,129){7}
//: {8}(273,184)(273,223){9}
//: {10}(275,225)(506,225)(506,272)(516,272){11}
//: {12}(271,225)(247,225){13}
wire w23;    //: /sn:0 /dp:1 {0}(460,104)(432,104){1}
wire w36;    //: /sn:0 {0}(207,179)(225,179){1}
wire w24;    //: /sn:0 {0}(127,174)(225,174){1}
wire w20;    //: /sn:0 {0}(246,99)(305,99)(305,98)(362,98){1}
wire w25;    //: /sn:0 /dp:1 {0}(295,150)(246,150){1}
wire w40;    //: /sn:0 /dp:1 {0}(516,277)(489,277){1}
wire w35;    //: /sn:0 /dp:1 {0}(468,279)(435,279){1}
wire w8;    //: /sn:0 {0}(127,224)(166,224)(166,222)(226,222){1}
wire w18;    //: /sn:0 {0}(161,300)(204,300)(204,301)(224,301){1}
wire w30;    //: /sn:0 {0}(203,101)(225,101){1}
wire w22;    //: /sn:0 /dp:1 {0}(411,101)(383,101){1}
wire w17;    //: /sn:0 {0}(127,296)(224,296){1}
wire w12;    //: /sn:0 {0}(161,254)(169,254)(169,253)(226,253){1}
wire w11;    //: /sn:0 {0}(127,246)(135,246)(135,248)(226,248){1}
wire w2;    //: /sn:0 {0}(127,96)(225,96){1}
wire w10;    //: /sn:0 {0}(161,152)(188,152){1}
wire w27;    //: /sn:0 /dp:1 {0}(347,180)(316,180){1}
wire w13;    //: /sn:0 {0}(247,251)(329,251){1}
//: {2}(333,251)(443,251)(443,274)(468,274){3}
//: {4}(331,249)(331,187){5}
//: {6}(333,185)(347,185){7}
//: {8}(331,183)(331,158)(346,158){9}
wire w33;    //: /sn:0 /dp:1 {0}(362,103)(345,103)(345,127)(316,127){1}
wire w5;    //: /sn:0 {0}(127,121)(225,121){1}
wire w29;    //: /sn:0 /dp:1 {0}(295,177)(246,177){1}
wire w9;    //: /sn:0 {0}(161,230)(169,230)(169,227)(226,227){1}
wire w39;    //: /sn:0 {0}(417,186)(450,186)(450,109)(460,109){1}
wire w26;    //: /sn:0 {0}(161,179)(191,179){1}
//: enddecls

  tran g8(.Z(w6), .I(B[2]));   //: @(155,126) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  tran g4(.Z(w2), .I(A[3]));   //: @(121,96) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  not g37 (.I(w26), .Z(w36));   //: @(197,179) /sn:0 /w:[ 1 0 ]
  not g34 (.I(w3), .Z(w30));   //: @(193,101) /sn:0 /w:[ 1 0 ]
  xnor g13 (.I0(w14), .I1(w15), .Z(w16));   //: @(236,276) /sn:0 /w:[ 1 1 0 ]
  and g3 (.I0(w2), .I1(w30), .Z(w20));   //: @(236,99) /sn:0 /w:[ 1 1 0 ]
  //: output g2 (AgB) @(604,107) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(86,76) /sn:0 /w:[ 0 ]
  tran g16(.Z(w12), .I(B[2]));   //: @(155,254) /sn:0 /R:2 /w:[ 0 12 11 ] /ss:1
  tran g11(.Z(w9), .I(B[3]));   //: @(155,230) /sn:0 /R:2 /w:[ 0 10 9 ] /ss:1
  and g28 (.I0(w29), .I1(w28), .Z(w27));   //: @(306,180) /sn:0 /w:[ 0 0 1 ]
  tran g10(.Z(w8), .I(A[3]));   //: @(121,224) /sn:0 /R:2 /w:[ 0 10 9 ] /ss:1
  tran g32(.Z(w24), .I(A[0]));   //: @(121,174) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  and g27 (.I0(w24), .I1(w36), .Z(w29));   //: @(236,177) /sn:0 /w:[ 1 1 1 ]
  tran g19(.Z(w17), .I(A[0]));   //: @(121,296) /sn:0 /R:2 /w:[ 0 16 15 ] /ss:1
  and g38 (.I0(w31), .I1(w16), .Z(w39));   //: @(407,186) /sn:0 /w:[ 0 5 0 ]
  and g6 (.I0(w5), .I1(w38), .Z(w4));   //: @(236,124) /sn:0 /w:[ 1 0 1 ]
  xnor g9 (.I0(w8), .I1(w9), .Z(w28));   //: @(237,225) /sn:0 /w:[ 1 1 13 ]
  tran g7(.Z(w5), .I(A[2]));   //: @(121,121) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  tran g31(.Z(w10), .I(B[1]));   //: @(155,152) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  tran g20(.Z(w18), .I(B[0]));   //: @(155,300) /sn:0 /R:2 /w:[ 0 16 15 ] /ss:1
  tran g15(.Z(w11), .I(A[2]));   //: @(121,246) /sn:0 /R:2 /w:[ 0 12 11 ] /ss:1
  //: joint g39 (w13) @(331, 185) /w:[ 6 8 -1 5 ]
  and g48 (.I0(w28), .I1(w40), .Z(AeqB));   //: @(527,275) /sn:0 /w:[ 11 0 1 ]
  //: output g43 (AeqB) @(611,275) /sn:0 /w:[ 0 ]
  //: joint g29 (w28) @(273, 182) /w:[ 1 2 -1 8 ]
  and g25 (.I0(w25), .I1(w28), .Z(w21));   //: @(306,153) /sn:0 /w:[ 0 5 1 ]
  tran g17(.Z(w14), .I(A[1]));   //: @(121,272) /sn:0 /R:2 /w:[ 0 14 13 ] /ss:1
  or g42 (.I0(w23), .I1(w39), .Z(AgB));   //: @(471,107) /sn:0 /w:[ 0 1 0 ]
  xnor g14 (.I0(w17), .I1(w18), .Z(w37));   //: @(235,299) /sn:0 /w:[ 1 1 1 ]
  tran g5(.Z(w3), .I(B[3]));   //: @(155,101) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: joint g47 (w13) @(331, 251) /w:[ 2 4 1 -1 ]
  and g44 (.I0(w16), .I1(w37), .Z(w35));   //: @(425,279) /sn:0 /w:[ 3 0 1 ]
  //: joint g21 (w28) @(273, 155) /w:[ 4 6 -1 3 ]
  not g36 (.I(w10), .Z(w34));   //: @(194,152) /sn:0 /w:[ 1 0 ]
  and g24 (.I0(w7), .I1(w34), .Z(w25));   //: @(236,150) /sn:0 /w:[ 1 1 1 ]
  or g41 (.I0(w22), .I1(w32), .Z(w23));   //: @(422,104) /sn:0 /w:[ 0 1 1 ]
  and g23 (.I0(w21), .I1(w13), .Z(w32));   //: @(357,156) /sn:0 /w:[ 0 9 0 ]
  or g40 (.I0(w20), .I1(w33), .Z(w22));   //: @(373,101) /sn:0 /w:[ 1 0 1 ]
  and g46 (.I0(w13), .I1(w35), .Z(w40));   //: @(479,277) /sn:0 /w:[ 3 0 1 ]
  //: joint g45 (w16) @(384, 276) /w:[ 2 4 1 -1 ]
  and g26 (.I0(w27), .I1(w13), .Z(w31));   //: @(358,183) /sn:0 /w:[ 0 7 1 ]
  not g35 (.I(w6), .Z(w38));   //: @(192,126) /sn:0 /w:[ 1 1 ]
  and g22 (.I0(w4), .I1(w28), .Z(w33));   //: @(306,127) /sn:0 /w:[ 0 7 1 ]
  //: input g0 (A) @(86,46) /sn:0 /w:[ 0 ]
  tran g18(.Z(w15), .I(B[1]));   //: @(155,278) /sn:0 /R:2 /w:[ 0 14 13 ] /ss:1
  xnor g12 (.I0(w11), .I1(w12), .Z(w13));   //: @(237,251) /sn:0 /w:[ 1 1 0 ]
  tran g33(.Z(w26), .I(B[0]));   //: @(155,179) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  tran g30(.Z(w7), .I(A[1]));   //: @(121,147) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  //: joint g49 (w28) @(273, 225) /w:[ 10 9 12 -1 ]

endmodule
